module AluDecoder
    (
    input logic alu_op, s,
    input logic [3:0] cmd,
    output logic no_write, shift,
    output logic [2:0] alu_ctl,
    output logic [1:0] flag_w
    );

    always_comb begin
        if (alu_op) begin
            case (cmd)
                4'b0100: {alu_ctl, no_write, shift} = 5'b000_0_0; // ADD
                4'b0010: {alu_ctl, no_write, shift} = 5'b001_0_0; // SUB
                4'b0000: {alu_ctl, no_write, shift} = 5'b010_0_0; // AND
                4'b1100: {alu_ctl, no_write, shift} = 5'b011_0_0; // OR
                4'b0101: {alu_ctl, no_write, shift} = 5'b100_0_0; // ADC
                4'b1010: {alu_ctl, no_write, shift} = 5'b001_1_0; // CMP
                4'b1011: {alu_ctl, no_write, shift} = 5'b000_1_0; // CMN
                4'b1000: {alu_ctl, no_write, shift} = 5'b010_1_0; // TST
                4'b1101: {alu_ctl, no_write, shift} = 5'b0xx_0_1; // LSL
                default: {alu_ctl, no_write, shift} = 5'bx; // not defined
            endcase

            flag_w[1] = s;
            flag_w[0] = s & (alu_ctl === 3'b000 | alu_ctl === 3'b001 | alu_ctl === 3'b100);
        end else begin
            alu_ctl = 3'b000;
            flag_w = 2'b00;
            no_write = 1'b0;
            shift = 1'b0;
        end
    end
endmodule
