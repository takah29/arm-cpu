module MainDecoder
    (
    input logic [1:0] op,
    input logic [5:0] funct,
    output logic branch, mem_to_reg, mem_w, alu_src, reg_w, alu_op, reg_src, post_idx,
    output logic [1:0] imm_src
    );

    logic [9:0] controls; // {branch, mem_to_reg, mem_w, alu_src, imm_src, reg_w, reg_src, alu_op, post_idx}

    function [9:0] dp_controls(input [5:0] funct);
        casex (funct)
            6'b0XXXXX: dp_controls = 10'b0_0_0_0_00_1_0_1_0; // DP Reg
            6'b1XXXXX: dp_controls = 10'b0_0_0_1_00_1_0_1_0; // DP Imm
            default: dp_controls = 10'bx;
        endcase
    endfunction

    function [9:0] mem_controls(input [5:0] funct);
        casex (funct)
            6'b01XX00: mem_controls = 10'b0_0_1_1_01_0_0_0_0; // STR (Imm)
            6'b11XX00: mem_controls = 10'b0_0_1_0_01_0_0_0_0; // STR (Reg)
            6'b01XX01: mem_controls = 10'b0_1_0_1_01_1_0_0_0; // LDR (Imm)
            6'b11XX01: mem_controls = 10'b0_1_0_0_01_1_0_0_0; // LDR (Reg)
            6'b00XX01: mem_controls = 10'b0_1_0_1_01_1_0_0_1; // LDR (Imm, PostIdx)
            6'b10XX01: mem_controls = 10'b0_1_0_0_01_1_0_0_1; // LDR (Reg, PostIdx)
            default: mem_controls = 10'bx;
        endcase
    endfunction

    always_comb begin
        case (op)
            2'b00: controls = dp_controls(funct); // DP
            2'b01: controls = mem_controls(funct); // Memory
            2'b10: controls = 10'b1_0_0_1_10_0_1_0_0; // B
            default: controls = 10'bx;
        endcase
    end

    assign {branch, mem_to_reg, mem_w, alu_src, imm_src, reg_w, reg_src, alu_op, post_idx} = controls;
endmodule
